typedef uvm_sequencer#(conter_transaction) counter_sequencer;