interface alu_if;
    logic[3:0] sig_if_s;
    logic[3:0] sig_if_a;
    logic[3:0] sig_if_b;
    logic sig_if_m;
    logic sig_if_c_in;
    logic[4:0] sig_if_f;
    logic clock;
endinterface