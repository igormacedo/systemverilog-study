module ram(
    data_in,
    data_out,
    addr,
    enable,
    read_write_en
);

input enable, read_write_en;


endmodule