module ramtb;