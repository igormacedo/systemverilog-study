interface counter_if;
    logic sig_if_clock;
    logic sig_if_reset;
    logic sig_if_clock_inhibit;
    logic sig_if_carry_out;
    logic[9:0] sig_if_number_bit;
endinterface