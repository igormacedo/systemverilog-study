typedef uvm_sequencer#(alu_transaction) alu_sequencer;