interface counter_if;
    logic sig_if_clock;
    logic sig_if_enable;
    logic[3:0] sig_if_value_in;
    logic[3:0] sig_if_out;
endinterface