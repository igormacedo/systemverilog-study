typedef uvm_sequencer#(counter_transaction) counter_sequencer;